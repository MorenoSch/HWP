-- analogToButtons
-- converts the reading of the adc into the corresponding button


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity analogToButtons is port(
	analogIn : in std_logic_vector(11 downto 0);
	
	Led: out std_logic_vector(5 downto 0)
);
end analogToButtons;


architecture behavior of analogToButtons is
begin
	-- TODO: add your code here
	
end behavior;